LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY MUX_CALCULATOR IS

	PORT (	SELECTOR  :    IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
				IN_1	    :	   IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
				IN_2	    :	   IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
				IN_3	    :	   IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
				OUTPUT    :	   OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
			
END ENTITY MUX_CALCULATOR;

ARCHITECTURE gateLevel OF MUX_CALCULATOR IS

				
BEGIN

	WITH SELECTOR SELECT
	
	OUTPUT <=  IN_1 WHEN "00",--MULTIPLICACION
				  IN_3 WHEN "01",--RESTA
				  IN_1 WHEN "10",--MULTIPLICACION
				  IN_2 WHEN "11";--SUMA

END ARCHITECTURE gateLevel;